// Verilog testbench created by TD v5.0.27252
// 2021-07-28 15:41:12

`timescale 1ns / 1ps

module TOP_tb();

reg CPLD_ATX_PWRGD;
reg CPLD_CASE_OPEN;
reg CPLD_CLK_25M;
reg CPLD_F_PANEL_PWRBTN;
reg CPLD_HW_RSTN;
reg CPLD_INT5_GPIO;
reg CPLD_INT6_GPIO;
reg CPLD_LPC_CLK_R;
reg CPLD_LPC_LFRAME;
reg CPLD_LPC_RST;
reg CPLD_SYS_WAKE_N;
reg CPLD_VDDQ_VPP_PG;
reg CPLD_VDD_CORE_P0V8_PG;
reg CPLD_VTT_PG;
reg FT_GPIO1_B3_CPLD;
reg FT_PWR_CTR0_CPLD;
reg FT_PWR_CTR1_CPLD;
wire CPLD_ALLMUTE_EC;
wire CPLD_BUZZER;
wire CPLD_FAN_PWM0;
wire CPLD_FAN_PWM1;
wire CPLD_FAN_PWM2;
wire CPLD_FAN_TACH0;
wire CPLD_FAN_TACH1;
wire CPLD_FAN_TACH2;
wire CPLD_FT_POR_N;
wire CPLD_FUSB_PWREN0;
wire CPLD_FUSB_PWREN1;
wire CPLD_GPIO_CASE0;
wire CPLD_GPIO_CASE1;
wire CPLD_HD_LED;
wire CPLD_LAN_PWR;
wire CPLD_MEM_RESET_S3;
wire CPLD_MUT_MONO_EC;
wire CPLD_P1V8_EN;
wire CPLD_PCIERST_SLOT;
wire CPLD_PCIE_LAN_RST_N;
wire CPLD_PWR_S0_EN;
wire CPLD_PWR_S3_EN;
wire CPLD_PWR_S4_S5_EN;
wire CPLD_RUSB_PWREN0;
wire CPLD_RUSB_PWREN1;
wire CPLD_SAFECARD_RSTN;
wire CPLD_SPKMUTE_EC;
wire CPLD_SYS_LED0;
wire CPLD_SYS_LED1;
wire CPLD_TCM_H_DISABLE;
wire CPLD_TCM_H_GPIO;
wire CPLD_TCM_H_PRESENT;
wire CPLD_TCM_ISORSTN;
wire CPLD_TCM_PORN;
wire CPLD_VDDQ_VPP_EN;
wire CPLD_VDD_CORE_EN;
wire CPLD_VTT_EN;
wire FT_GPIO0_A1;
wire HD_LED_FP;
wire SYS_S3N_CPLD;
wire SYS_S5N_CPLD;
wire CPLD_CLKGEN_CLK;
wire CPLD_CLKGEN_DAT;
wire CPLD_I2C1_SCL;
wire CPLD_I2C1_SDA;
wire CPLD_LPC_IRQ;
wire [3:0] CPLD_LPC_LAD;
wire CPLD_SCL_TEMP;
wire CPLD_SDA_TEMP;
wire CPLD_SLOT_I2C_CLK;
wire CPLD_SLOT_I2C_SDA;
wire SCI_CPLD;

//Clock process
parameter PERIOD = 10;
always #(PERIOD/2) CPLD_SLOT_I2C_CLK = ~CPLD_SLOT_I2C_CLK;

//glbl Instantiate
glbl glbl();

//Unit Instantiate
TOP uut(
	.CPLD_ATX_PWRGD(CPLD_ATX_PWRGD),
	.CPLD_CASE_OPEN(CPLD_CASE_OPEN),
	.CPLD_CLK_25M(CPLD_CLK_25M),
	.CPLD_F_PANEL_PWRBTN(CPLD_F_PANEL_PWRBTN),
	.CPLD_HW_RSTN(CPLD_HW_RSTN),
	.CPLD_INT5_GPIO(CPLD_INT5_GPIO),
	.CPLD_INT6_GPIO(CPLD_INT6_GPIO),
	.CPLD_LPC_CLK_R(CPLD_LPC_CLK_R),
	.CPLD_LPC_LFRAME(CPLD_LPC_LFRAME),
	.CPLD_LPC_RST(CPLD_LPC_RST),
	.CPLD_SYS_WAKE_N(CPLD_SYS_WAKE_N),
	.CPLD_VDDQ_VPP_PG(CPLD_VDDQ_VPP_PG),
	.CPLD_VDD_CORE_P0V8_PG(CPLD_VDD_CORE_P0V8_PG),
	.CPLD_VTT_PG(CPLD_VTT_PG),
	.FT_GPIO1_B3_CPLD(FT_GPIO1_B3_CPLD),
	.FT_PWR_CTR0_CPLD(FT_PWR_CTR0_CPLD),
	.FT_PWR_CTR1_CPLD(FT_PWR_CTR1_CPLD),
	.CPLD_ALLMUTE_EC(CPLD_ALLMUTE_EC),
	.CPLD_BUZZER(CPLD_BUZZER),
	.CPLD_FAN_PWM0(CPLD_FAN_PWM0),
	.CPLD_FAN_PWM1(CPLD_FAN_PWM1),
	.CPLD_FAN_PWM2(CPLD_FAN_PWM2),
	.CPLD_FAN_TACH0(CPLD_FAN_TACH0),
	.CPLD_FAN_TACH1(CPLD_FAN_TACH1),
	.CPLD_FAN_TACH2(CPLD_FAN_TACH2),
	.CPLD_FT_POR_N(CPLD_FT_POR_N),
	.CPLD_FUSB_PWREN0(CPLD_FUSB_PWREN0),
	.CPLD_FUSB_PWREN1(CPLD_FUSB_PWREN1),
	.CPLD_GPIO_CASE0(CPLD_GPIO_CASE0),
	.CPLD_GPIO_CASE1(CPLD_GPIO_CASE1),
	.CPLD_HD_LED(CPLD_HD_LED),
	.CPLD_LAN_PWR(CPLD_LAN_PWR),
	.CPLD_MEM_RESET_S3(CPLD_MEM_RESET_S3),
	.CPLD_MUT_MONO_EC(CPLD_MUT_MONO_EC),
	.CPLD_P1V8_EN(CPLD_P1V8_EN),
	.CPLD_PCIERST_SLOT(CPLD_PCIERST_SLOT),
	.CPLD_PCIE_LAN_RST_N(CPLD_PCIE_LAN_RST_N),
	.CPLD_PWR_S0_EN(CPLD_PWR_S0_EN),
	.CPLD_PWR_S3_EN(CPLD_PWR_S3_EN),
	.CPLD_PWR_S4_S5_EN(CPLD_PWR_S4_S5_EN),
	.CPLD_RUSB_PWREN0(CPLD_RUSB_PWREN0),
	.CPLD_RUSB_PWREN1(CPLD_RUSB_PWREN1),
	.CPLD_SAFECARD_RSTN(CPLD_SAFECARD_RSTN),
	.CPLD_SPKMUTE_EC(CPLD_SPKMUTE_EC),
	.CPLD_SYS_LED0(CPLD_SYS_LED0),
	.CPLD_SYS_LED1(CPLD_SYS_LED1),
	.CPLD_TCM_H_DISABLE(CPLD_TCM_H_DISABLE),
	.CPLD_TCM_H_GPIO(CPLD_TCM_H_GPIO),
	.CPLD_TCM_H_PRESENT(CPLD_TCM_H_PRESENT),
	.CPLD_TCM_ISORSTN(CPLD_TCM_ISORSTN),
	.CPLD_TCM_PORN(CPLD_TCM_PORN),
	.CPLD_VDDQ_VPP_EN(CPLD_VDDQ_VPP_EN),
	.CPLD_VDD_CORE_EN(CPLD_VDD_CORE_EN),
	.CPLD_VTT_EN(CPLD_VTT_EN),
	.FT_GPIO0_A1(FT_GPIO0_A1),
	.HD_LED_FP(HD_LED_FP),
	.SYS_S3N_CPLD(SYS_S3N_CPLD),
	.SYS_S5N_CPLD(SYS_S5N_CPLD),
	.CPLD_CLKGEN_CLK(CPLD_CLKGEN_CLK),
	.CPLD_CLKGEN_DAT(CPLD_CLKGEN_DAT),
	.CPLD_I2C1_SCL(CPLD_I2C1_SCL),
	.CPLD_I2C1_SDA(CPLD_I2C1_SDA),
	.CPLD_LPC_IRQ(CPLD_LPC_IRQ),
	.CPLD_LPC_LAD(CPLD_LPC_LAD),
	.CPLD_SCL_TEMP(CPLD_SCL_TEMP),
	.CPLD_SDA_TEMP(CPLD_SDA_TEMP),
	.CPLD_SLOT_I2C_CLK(CPLD_SLOT_I2C_CLK),
	.CPLD_SLOT_I2C_SDA(CPLD_SLOT_I2C_SDA),
	.SCI_CPLD(SCI_CPLD));

//Stimulus process
initial begin
//To be inserted
end

endmodule